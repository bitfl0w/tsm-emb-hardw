-- lab3_sopc.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity lab3_sopc is
	port (
		buttons_export        : inout std_logic_vector(7 downto 0)  := (others => '0'); --         buttons.export
		clk_clk               : in    std_logic                     := '0';             --             clk.clk
		led_row2_export       : inout std_logic_vector(7 downto 0)  := (others => '0'); --        led_row2.export
		led_row3_export       : inout std_logic_vector(7 downto 0)  := (others => '0'); --        led_row3.export
		reset_reset_n         : in    std_logic                     := '0';             --           reset.reset_n
		sdram_clk_clk         : out   std_logic;                                        --       sdram_clk.clk
		sdram_ctrl_wire_addr  : out   std_logic_vector(11 downto 0);                    -- sdram_ctrl_wire.addr
		sdram_ctrl_wire_ba    : out   std_logic_vector(1 downto 0);                     --                .ba
		sdram_ctrl_wire_cas_n : out   std_logic;                                        --                .cas_n
		sdram_ctrl_wire_cke   : out   std_logic;                                        --                .cke
		sdram_ctrl_wire_cs_n  : out   std_logic;                                        --                .cs_n
		sdram_ctrl_wire_dq    : inout std_logic_vector(15 downto 0) := (others => '0'); --                .dq
		sdram_ctrl_wire_dqm   : out   std_logic_vector(1 downto 0);                     --                .dqm
		sdram_ctrl_wire_ras_n : out   std_logic;                                        --                .ras_n
		sdram_ctrl_wire_we_n  : out   std_logic                                         --                .we_n
	);
end entity lab3_sopc;

architecture rtl of lab3_sopc is
	component lab3_sopc_CPU is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(25 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(25 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component lab3_sopc_CPU;

	component lab3_sopc_PLL is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c2                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component lab3_sopc_PLL;

	component lab3_sopc_SDRAM_ctrl is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(22 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component lab3_sopc_SDRAM_ctrl;

	component lab3_sopc_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component lab3_sopc_jtag_uart;

	component simplePIO is
		port (
			irq          : out   std_logic;                                       -- irq
			av_address   : in    std_logic_vector(2 downto 0) := (others => 'X'); -- address
			av_read      : in    std_logic                    := 'X';             -- read
			av_readdata  : out   std_logic_vector(7 downto 0);                    -- readdata
			av_write     : in    std_logic                    := 'X';             -- write
			av_writedata : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			conduit_data : inout std_logic_vector(7 downto 0) := (others => 'X'); -- export
			clk          : in    std_logic                    := 'X';             -- clk
			reset_n      : in    std_logic                    := 'X'              -- reset_n
		);
	end component simplePIO;

	component lab3_sopc_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component lab3_sopc_sysid;

	component lab3_sopc_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                           : in  std_logic                     := 'X';             -- clk
			PLL_c0_clk                                              : in  std_logic                     := 'X';             -- clk
			CPU_reset_reset_bridge_in_reset_reset                   : in  std_logic                     := 'X';             -- reset
			jtag_uart_reset_reset_bridge_in_reset_reset             : in  std_logic                     := 'X';             -- reset
			parallel_port_buttons_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			PLL_inclk_interface_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			CPU_data_master_address                                 : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			CPU_data_master_waitrequest                             : out std_logic;                                        -- waitrequest
			CPU_data_master_byteenable                              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			CPU_data_master_read                                    : in  std_logic                     := 'X';             -- read
			CPU_data_master_readdata                                : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_data_master_readdatavalid                           : out std_logic;                                        -- readdatavalid
			CPU_data_master_write                                   : in  std_logic                     := 'X';             -- write
			CPU_data_master_writedata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			CPU_data_master_debugaccess                             : in  std_logic                     := 'X';             -- debugaccess
			CPU_instruction_master_address                          : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			CPU_instruction_master_waitrequest                      : out std_logic;                                        -- waitrequest
			CPU_instruction_master_read                             : in  std_logic                     := 'X';             -- read
			CPU_instruction_master_readdata                         : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_instruction_master_readdatavalid                    : out std_logic;                                        -- readdatavalid
			CPU_debug_mem_slave_address                             : out std_logic_vector(8 downto 0);                     -- address
			CPU_debug_mem_slave_write                               : out std_logic;                                        -- write
			CPU_debug_mem_slave_read                                : out std_logic;                                        -- read
			CPU_debug_mem_slave_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			CPU_debug_mem_slave_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			CPU_debug_mem_slave_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			CPU_debug_mem_slave_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			CPU_debug_mem_slave_debugaccess                         : out std_logic;                                        -- debugaccess
			jtag_uart_avalon_jtag_slave_address                     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                       : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                        : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest                 : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                  : out std_logic;                                        -- chipselect
			parallel_port_buttons_av_address                        : out std_logic_vector(2 downto 0);                     -- address
			parallel_port_buttons_av_write                          : out std_logic;                                        -- write
			parallel_port_buttons_av_read                           : out std_logic;                                        -- read
			parallel_port_buttons_av_readdata                       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			parallel_port_buttons_av_writedata                      : out std_logic_vector(7 downto 0);                     -- writedata
			parallel_port_led_row2_av_address                       : out std_logic_vector(2 downto 0);                     -- address
			parallel_port_led_row2_av_write                         : out std_logic;                                        -- write
			parallel_port_led_row2_av_read                          : out std_logic;                                        -- read
			parallel_port_led_row2_av_readdata                      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			parallel_port_led_row2_av_writedata                     : out std_logic_vector(7 downto 0);                     -- writedata
			parallel_port_led_row3_av_address                       : out std_logic_vector(2 downto 0);                     -- address
			parallel_port_led_row3_av_write                         : out std_logic;                                        -- write
			parallel_port_led_row3_av_read                          : out std_logic;                                        -- read
			parallel_port_led_row3_av_readdata                      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			parallel_port_led_row3_av_writedata                     : out std_logic_vector(7 downto 0);                     -- writedata
			PLL_pll_slave_address                                   : out std_logic_vector(1 downto 0);                     -- address
			PLL_pll_slave_write                                     : out std_logic;                                        -- write
			PLL_pll_slave_read                                      : out std_logic;                                        -- read
			PLL_pll_slave_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PLL_pll_slave_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			SDRAM_ctrl_s1_address                                   : out std_logic_vector(22 downto 0);                    -- address
			SDRAM_ctrl_s1_write                                     : out std_logic;                                        -- write
			SDRAM_ctrl_s1_read                                      : out std_logic;                                        -- read
			SDRAM_ctrl_s1_readdata                                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SDRAM_ctrl_s1_writedata                                 : out std_logic_vector(15 downto 0);                    -- writedata
			SDRAM_ctrl_s1_byteenable                                : out std_logic_vector(1 downto 0);                     -- byteenable
			SDRAM_ctrl_s1_readdatavalid                             : in  std_logic                     := 'X';             -- readdatavalid
			SDRAM_ctrl_s1_waitrequest                               : in  std_logic                     := 'X';             -- waitrequest
			SDRAM_ctrl_s1_chipselect                                : out std_logic;                                        -- chipselect
			sysid_control_slave_address                             : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component lab3_sopc_mm_interconnect_0;

	component lab3_sopc_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component lab3_sopc_irq_mapper;

	component lab3_sopc_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component lab3_sopc_rst_controller;

	component lab3_sopc_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component lab3_sopc_rst_controller_001;

	component lab3_sopc_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component lab3_sopc_rst_controller_002;

	signal pll_c0_clk                                                    : std_logic;                     -- PLL:c0 -> [CPU:clk, SDRAM_ctrl:clk, irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:PLL_c0_clk, parallel_port_buttons:clk, parallel_port_led_row2:clk, parallel_port_led_row3:clk, rst_controller:clk, rst_controller_002:clk, sysid:clock]
	signal cpu_debug_reset_request_reset                                 : std_logic;                     -- CPU:debug_reset_request -> [cpu_debug_reset_request_reset:in, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal cpu_data_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	signal cpu_data_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	signal cpu_data_master_debugaccess                                   : std_logic;                     -- CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	signal cpu_data_master_address                                       : std_logic_vector(25 downto 0); -- CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	signal cpu_data_master_byteenable                                    : std_logic_vector(3 downto 0);  -- CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	signal cpu_data_master_read                                          : std_logic;                     -- CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	signal cpu_data_master_readdatavalid                                 : std_logic;                     -- mm_interconnect_0:CPU_data_master_readdatavalid -> CPU:d_readdatavalid
	signal cpu_data_master_write                                         : std_logic;                     -- CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	signal cpu_data_master_writedata                                     : std_logic_vector(31 downto 0); -- CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	signal cpu_instruction_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	signal cpu_instruction_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	signal cpu_instruction_master_address                                : std_logic_vector(25 downto 0); -- CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	signal cpu_instruction_master_read                                   : std_logic;                     -- CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	signal cpu_instruction_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:CPU_instruction_master_readdatavalid -> CPU:i_readdatavalid
	signal mm_interconnect_0_parallel_port_buttons_av_readdata           : std_logic_vector(7 downto 0);  -- parallel_port_buttons:av_readdata -> mm_interconnect_0:parallel_port_buttons_av_readdata
	signal mm_interconnect_0_parallel_port_buttons_av_address            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:parallel_port_buttons_av_address -> parallel_port_buttons:av_address
	signal mm_interconnect_0_parallel_port_buttons_av_read               : std_logic;                     -- mm_interconnect_0:parallel_port_buttons_av_read -> parallel_port_buttons:av_read
	signal mm_interconnect_0_parallel_port_buttons_av_write              : std_logic;                     -- mm_interconnect_0:parallel_port_buttons_av_write -> parallel_port_buttons:av_write
	signal mm_interconnect_0_parallel_port_buttons_av_writedata          : std_logic_vector(7 downto 0);  -- mm_interconnect_0:parallel_port_buttons_av_writedata -> parallel_port_buttons:av_writedata
	signal mm_interconnect_0_parallel_port_led_row2_av_readdata          : std_logic_vector(7 downto 0);  -- parallel_port_led_row2:av_readdata -> mm_interconnect_0:parallel_port_led_row2_av_readdata
	signal mm_interconnect_0_parallel_port_led_row2_av_address           : std_logic_vector(2 downto 0);  -- mm_interconnect_0:parallel_port_led_row2_av_address -> parallel_port_led_row2:av_address
	signal mm_interconnect_0_parallel_port_led_row2_av_read              : std_logic;                     -- mm_interconnect_0:parallel_port_led_row2_av_read -> parallel_port_led_row2:av_read
	signal mm_interconnect_0_parallel_port_led_row2_av_write             : std_logic;                     -- mm_interconnect_0:parallel_port_led_row2_av_write -> parallel_port_led_row2:av_write
	signal mm_interconnect_0_parallel_port_led_row2_av_writedata         : std_logic_vector(7 downto 0);  -- mm_interconnect_0:parallel_port_led_row2_av_writedata -> parallel_port_led_row2:av_writedata
	signal mm_interconnect_0_parallel_port_led_row3_av_readdata          : std_logic_vector(7 downto 0);  -- parallel_port_led_row3:av_readdata -> mm_interconnect_0:parallel_port_led_row3_av_readdata
	signal mm_interconnect_0_parallel_port_led_row3_av_address           : std_logic_vector(2 downto 0);  -- mm_interconnect_0:parallel_port_led_row3_av_address -> parallel_port_led_row3:av_address
	signal mm_interconnect_0_parallel_port_led_row3_av_read              : std_logic;                     -- mm_interconnect_0:parallel_port_led_row3_av_read -> parallel_port_led_row3:av_read
	signal mm_interconnect_0_parallel_port_led_row3_av_write             : std_logic;                     -- mm_interconnect_0:parallel_port_led_row3_av_write -> parallel_port_led_row3:av_write
	signal mm_interconnect_0_parallel_port_led_row3_av_writedata         : std_logic_vector(7 downto 0);  -- mm_interconnect_0:parallel_port_led_row3_av_writedata -> parallel_port_led_row3:av_writedata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_sysid_control_slave_readdata                : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                 : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                : std_logic_vector(31 downto 0); -- CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest             : std_logic;                     -- CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess             : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                 : std_logic_vector(8 downto 0);  -- mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                    : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                   : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	signal mm_interconnect_0_pll_pll_slave_readdata                      : std_logic_vector(31 downto 0); -- PLL:readdata -> mm_interconnect_0:PLL_pll_slave_readdata
	signal mm_interconnect_0_pll_pll_slave_address                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:PLL_pll_slave_address -> PLL:address
	signal mm_interconnect_0_pll_pll_slave_read                          : std_logic;                     -- mm_interconnect_0:PLL_pll_slave_read -> PLL:read
	signal mm_interconnect_0_pll_pll_slave_write                         : std_logic;                     -- mm_interconnect_0:PLL_pll_slave_write -> PLL:write
	signal mm_interconnect_0_pll_pll_slave_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:PLL_pll_slave_writedata -> PLL:writedata
	signal mm_interconnect_0_sdram_ctrl_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:SDRAM_ctrl_s1_chipselect -> SDRAM_ctrl:az_cs
	signal mm_interconnect_0_sdram_ctrl_s1_readdata                      : std_logic_vector(15 downto 0); -- SDRAM_ctrl:za_data -> mm_interconnect_0:SDRAM_ctrl_s1_readdata
	signal mm_interconnect_0_sdram_ctrl_s1_waitrequest                   : std_logic;                     -- SDRAM_ctrl:za_waitrequest -> mm_interconnect_0:SDRAM_ctrl_s1_waitrequest
	signal mm_interconnect_0_sdram_ctrl_s1_address                       : std_logic_vector(22 downto 0); -- mm_interconnect_0:SDRAM_ctrl_s1_address -> SDRAM_ctrl:az_addr
	signal mm_interconnect_0_sdram_ctrl_s1_read                          : std_logic;                     -- mm_interconnect_0:SDRAM_ctrl_s1_read -> mm_interconnect_0_sdram_ctrl_s1_read:in
	signal mm_interconnect_0_sdram_ctrl_s1_byteenable                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SDRAM_ctrl_s1_byteenable -> mm_interconnect_0_sdram_ctrl_s1_byteenable:in
	signal mm_interconnect_0_sdram_ctrl_s1_readdatavalid                 : std_logic;                     -- SDRAM_ctrl:za_valid -> mm_interconnect_0:SDRAM_ctrl_s1_readdatavalid
	signal mm_interconnect_0_sdram_ctrl_s1_write                         : std_logic;                     -- mm_interconnect_0:SDRAM_ctrl_s1_write -> mm_interconnect_0_sdram_ctrl_s1_write:in
	signal mm_interconnect_0_sdram_ctrl_s1_writedata                     : std_logic_vector(15 downto 0); -- mm_interconnect_0:SDRAM_ctrl_s1_writedata -> SDRAM_ctrl:az_data
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- parallel_port_buttons:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- parallel_port_led_row2:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                      : std_logic;                     -- parallel_port_led_row3:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver3_irq
	signal cpu_irq_irq                                                   : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> CPU:irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [CPU:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                            : std_logic;                     -- rst_controller_001:reset_out -> [PLL:reset, mm_interconnect_0:PLL_inclk_interface_reset_reset_bridge_in_reset_reset]
	signal rst_controller_002_reset_out_reset                            : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:parallel_port_buttons_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in]
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal cpu_debug_reset_request_reset_ports_inv                       : std_logic;                     -- cpu_debug_reset_request_reset:inv -> jtag_uart:rst_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_sdram_ctrl_s1_read_ports_inv                : std_logic;                     -- mm_interconnect_0_sdram_ctrl_s1_read:inv -> SDRAM_ctrl:az_rd_n
	signal mm_interconnect_0_sdram_ctrl_s1_byteenable_ports_inv          : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_ctrl_s1_byteenable:inv -> SDRAM_ctrl:az_be_n
	signal mm_interconnect_0_sdram_ctrl_s1_write_ports_inv               : std_logic;                     -- mm_interconnect_0_sdram_ctrl_s1_write:inv -> SDRAM_ctrl:az_wr_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [CPU:reset_n, SDRAM_ctrl:reset_n, sysid:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> [parallel_port_buttons:reset_n, parallel_port_led_row2:reset_n, parallel_port_led_row3:reset_n]

begin

	cpu : component lab3_sopc_CPU
		port map (
			clk                                 => pll_c0_clk,                                        --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	pll : component lab3_sopc_PLL
		port map (
			clk                => clk_clk,                                   --       inclk_interface.clk
			reset              => rst_controller_001_reset_out_reset,        -- inclk_interface_reset.reset
			read               => mm_interconnect_0_pll_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_pll_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_pll_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_pll_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_pll_pll_slave_writedata, --                      .writedata
			c0                 => pll_c0_clk,                                --                    c0.clk
			c2                 => sdram_clk_clk,                             --                    c2.clk
			scandone           => open,                                      --           (terminated)
			scandataout        => open,                                      --           (terminated)
			areset             => '0',                                       --           (terminated)
			locked             => open,                                      --           (terminated)
			phasedone          => open,                                      --           (terminated)
			phasecounterselect => "0000",                                    --           (terminated)
			phaseupdown        => '0',                                       --           (terminated)
			phasestep          => '0',                                       --           (terminated)
			scanclk            => '0',                                       --           (terminated)
			scanclkena         => '0',                                       --           (terminated)
			scandata           => '0',                                       --           (terminated)
			configupdate       => '0'                                        --           (terminated)
		);

	sdram_ctrl : component lab3_sopc_SDRAM_ctrl
		port map (
			clk            => pll_c0_clk,                                           --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,             -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_ctrl_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_ctrl_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_ctrl_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_ctrl_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_ctrl_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_ctrl_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_ctrl_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_ctrl_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_ctrl_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_ctrl_wire_addr,                                 --  wire.export
			zs_ba          => sdram_ctrl_wire_ba,                                   --      .export
			zs_cas_n       => sdram_ctrl_wire_cas_n,                                --      .export
			zs_cke         => sdram_ctrl_wire_cke,                                  --      .export
			zs_cs_n        => sdram_ctrl_wire_cs_n,                                 --      .export
			zs_dq          => sdram_ctrl_wire_dq,                                   --      .export
			zs_dqm         => sdram_ctrl_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_ctrl_wire_ras_n,                                --      .export
			zs_we_n        => sdram_ctrl_wire_we_n                                  --      .export
		);

	jtag_uart : component lab3_sopc_jtag_uart
		port map (
			clk            => pll_c0_clk,                                                    --               clk.clk
			rst_n          => cpu_debug_reset_request_reset_ports_inv,                       --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver3_irq                                       --               irq.irq
		);

	parallel_port_buttons : component simplePIO
		port map (
			irq          => irq_mapper_receiver0_irq,                             -- interrupt_sender.irq
			av_address   => mm_interconnect_0_parallel_port_buttons_av_address,   --               av.address
			av_read      => mm_interconnect_0_parallel_port_buttons_av_read,      --                 .read
			av_readdata  => mm_interconnect_0_parallel_port_buttons_av_readdata,  --                 .readdata
			av_write     => mm_interconnect_0_parallel_port_buttons_av_write,     --                 .write
			av_writedata => mm_interconnect_0_parallel_port_buttons_av_writedata, --                 .writedata
			conduit_data => buttons_export,                                       --         pio_port.export
			clk          => pll_c0_clk,                                           --            clock.clk
			reset_n      => rst_controller_002_reset_out_reset_ports_inv          --            reset.reset_n
		);

	parallel_port_led_row2 : component simplePIO
		port map (
			irq          => irq_mapper_receiver1_irq,                              -- interrupt_sender.irq
			av_address   => mm_interconnect_0_parallel_port_led_row2_av_address,   --               av.address
			av_read      => mm_interconnect_0_parallel_port_led_row2_av_read,      --                 .read
			av_readdata  => mm_interconnect_0_parallel_port_led_row2_av_readdata,  --                 .readdata
			av_write     => mm_interconnect_0_parallel_port_led_row2_av_write,     --                 .write
			av_writedata => mm_interconnect_0_parallel_port_led_row2_av_writedata, --                 .writedata
			conduit_data => led_row2_export,                                       --         pio_port.export
			clk          => pll_c0_clk,                                            --            clock.clk
			reset_n      => rst_controller_002_reset_out_reset_ports_inv           --            reset.reset_n
		);

	parallel_port_led_row3 : component simplePIO
		port map (
			irq          => irq_mapper_receiver2_irq,                              -- interrupt_sender.irq
			av_address   => mm_interconnect_0_parallel_port_led_row3_av_address,   --               av.address
			av_read      => mm_interconnect_0_parallel_port_led_row3_av_read,      --                 .read
			av_readdata  => mm_interconnect_0_parallel_port_led_row3_av_readdata,  --                 .readdata
			av_write     => mm_interconnect_0_parallel_port_led_row3_av_write,     --                 .write
			av_writedata => mm_interconnect_0_parallel_port_led_row3_av_writedata, --                 .writedata
			conduit_data => led_row3_export,                                       --         pio_port.export
			clk          => pll_c0_clk,                                            --            clock.clk
			reset_n      => rst_controller_002_reset_out_reset_ports_inv           --            reset.reset_n
		);

	sysid : component lab3_sopc_sysid
		port map (
			clock    => pll_c0_clk,                                       --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component lab3_sopc_mm_interconnect_0
		port map (
			clk_0_clk_clk                                           => clk_clk,                                                   --                                         clk_0_clk.clk
			PLL_c0_clk                                              => pll_c0_clk,                                                --                                            PLL_c0.clk
			CPU_reset_reset_bridge_in_reset_reset                   => rst_controller_reset_out_reset,                            --                   CPU_reset_reset_bridge_in_reset.reset
			jtag_uart_reset_reset_bridge_in_reset_reset             => cpu_debug_reset_request_reset,                             --             jtag_uart_reset_reset_bridge_in_reset.reset
			parallel_port_buttons_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                        -- parallel_port_buttons_reset_reset_bridge_in_reset.reset
			PLL_inclk_interface_reset_reset_bridge_in_reset_reset   => rst_controller_001_reset_out_reset,                        --   PLL_inclk_interface_reset_reset_bridge_in_reset.reset
			CPU_data_master_address                                 => cpu_data_master_address,                                   --                                   CPU_data_master.address
			CPU_data_master_waitrequest                             => cpu_data_master_waitrequest,                               --                                                  .waitrequest
			CPU_data_master_byteenable                              => cpu_data_master_byteenable,                                --                                                  .byteenable
			CPU_data_master_read                                    => cpu_data_master_read,                                      --                                                  .read
			CPU_data_master_readdata                                => cpu_data_master_readdata,                                  --                                                  .readdata
			CPU_data_master_readdatavalid                           => cpu_data_master_readdatavalid,                             --                                                  .readdatavalid
			CPU_data_master_write                                   => cpu_data_master_write,                                     --                                                  .write
			CPU_data_master_writedata                               => cpu_data_master_writedata,                                 --                                                  .writedata
			CPU_data_master_debugaccess                             => cpu_data_master_debugaccess,                               --                                                  .debugaccess
			CPU_instruction_master_address                          => cpu_instruction_master_address,                            --                            CPU_instruction_master.address
			CPU_instruction_master_waitrequest                      => cpu_instruction_master_waitrequest,                        --                                                  .waitrequest
			CPU_instruction_master_read                             => cpu_instruction_master_read,                               --                                                  .read
			CPU_instruction_master_readdata                         => cpu_instruction_master_readdata,                           --                                                  .readdata
			CPU_instruction_master_readdatavalid                    => cpu_instruction_master_readdatavalid,                      --                                                  .readdatavalid
			CPU_debug_mem_slave_address                             => mm_interconnect_0_cpu_debug_mem_slave_address,             --                               CPU_debug_mem_slave.address
			CPU_debug_mem_slave_write                               => mm_interconnect_0_cpu_debug_mem_slave_write,               --                                                  .write
			CPU_debug_mem_slave_read                                => mm_interconnect_0_cpu_debug_mem_slave_read,                --                                                  .read
			CPU_debug_mem_slave_readdata                            => mm_interconnect_0_cpu_debug_mem_slave_readdata,            --                                                  .readdata
			CPU_debug_mem_slave_writedata                           => mm_interconnect_0_cpu_debug_mem_slave_writedata,           --                                                  .writedata
			CPU_debug_mem_slave_byteenable                          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,          --                                                  .byteenable
			CPU_debug_mem_slave_waitrequest                         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,         --                                                  .waitrequest
			CPU_debug_mem_slave_debugaccess                         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,         --                                                  .debugaccess
			jtag_uart_avalon_jtag_slave_address                     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --                       jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                                  .write
			jtag_uart_avalon_jtag_slave_read                        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                                  .read
			jtag_uart_avalon_jtag_slave_readdata                    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                                  .readdata
			jtag_uart_avalon_jtag_slave_writedata                   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                                  .writedata
			jtag_uart_avalon_jtag_slave_waitrequest                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                                  .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                                  .chipselect
			parallel_port_buttons_av_address                        => mm_interconnect_0_parallel_port_buttons_av_address,        --                          parallel_port_buttons_av.address
			parallel_port_buttons_av_write                          => mm_interconnect_0_parallel_port_buttons_av_write,          --                                                  .write
			parallel_port_buttons_av_read                           => mm_interconnect_0_parallel_port_buttons_av_read,           --                                                  .read
			parallel_port_buttons_av_readdata                       => mm_interconnect_0_parallel_port_buttons_av_readdata,       --                                                  .readdata
			parallel_port_buttons_av_writedata                      => mm_interconnect_0_parallel_port_buttons_av_writedata,      --                                                  .writedata
			parallel_port_led_row2_av_address                       => mm_interconnect_0_parallel_port_led_row2_av_address,       --                         parallel_port_led_row2_av.address
			parallel_port_led_row2_av_write                         => mm_interconnect_0_parallel_port_led_row2_av_write,         --                                                  .write
			parallel_port_led_row2_av_read                          => mm_interconnect_0_parallel_port_led_row2_av_read,          --                                                  .read
			parallel_port_led_row2_av_readdata                      => mm_interconnect_0_parallel_port_led_row2_av_readdata,      --                                                  .readdata
			parallel_port_led_row2_av_writedata                     => mm_interconnect_0_parallel_port_led_row2_av_writedata,     --                                                  .writedata
			parallel_port_led_row3_av_address                       => mm_interconnect_0_parallel_port_led_row3_av_address,       --                         parallel_port_led_row3_av.address
			parallel_port_led_row3_av_write                         => mm_interconnect_0_parallel_port_led_row3_av_write,         --                                                  .write
			parallel_port_led_row3_av_read                          => mm_interconnect_0_parallel_port_led_row3_av_read,          --                                                  .read
			parallel_port_led_row3_av_readdata                      => mm_interconnect_0_parallel_port_led_row3_av_readdata,      --                                                  .readdata
			parallel_port_led_row3_av_writedata                     => mm_interconnect_0_parallel_port_led_row3_av_writedata,     --                                                  .writedata
			PLL_pll_slave_address                                   => mm_interconnect_0_pll_pll_slave_address,                   --                                     PLL_pll_slave.address
			PLL_pll_slave_write                                     => mm_interconnect_0_pll_pll_slave_write,                     --                                                  .write
			PLL_pll_slave_read                                      => mm_interconnect_0_pll_pll_slave_read,                      --                                                  .read
			PLL_pll_slave_readdata                                  => mm_interconnect_0_pll_pll_slave_readdata,                  --                                                  .readdata
			PLL_pll_slave_writedata                                 => mm_interconnect_0_pll_pll_slave_writedata,                 --                                                  .writedata
			SDRAM_ctrl_s1_address                                   => mm_interconnect_0_sdram_ctrl_s1_address,                   --                                     SDRAM_ctrl_s1.address
			SDRAM_ctrl_s1_write                                     => mm_interconnect_0_sdram_ctrl_s1_write,                     --                                                  .write
			SDRAM_ctrl_s1_read                                      => mm_interconnect_0_sdram_ctrl_s1_read,                      --                                                  .read
			SDRAM_ctrl_s1_readdata                                  => mm_interconnect_0_sdram_ctrl_s1_readdata,                  --                                                  .readdata
			SDRAM_ctrl_s1_writedata                                 => mm_interconnect_0_sdram_ctrl_s1_writedata,                 --                                                  .writedata
			SDRAM_ctrl_s1_byteenable                                => mm_interconnect_0_sdram_ctrl_s1_byteenable,                --                                                  .byteenable
			SDRAM_ctrl_s1_readdatavalid                             => mm_interconnect_0_sdram_ctrl_s1_readdatavalid,             --                                                  .readdatavalid
			SDRAM_ctrl_s1_waitrequest                               => mm_interconnect_0_sdram_ctrl_s1_waitrequest,               --                                                  .waitrequest
			SDRAM_ctrl_s1_chipselect                                => mm_interconnect_0_sdram_ctrl_s1_chipselect,                --                                                  .chipselect
			sysid_control_slave_address                             => mm_interconnect_0_sysid_control_slave_address,             --                               sysid_control_slave.address
			sysid_control_slave_readdata                            => mm_interconnect_0_sysid_control_slave_readdata             --                                                  .readdata
		);

	irq_mapper : component lab3_sopc_irq_mapper
		port map (
			clk           => pll_c0_clk,                     --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			sender_irq    => cpu_irq_irq                     --    sender.irq
		);

	rst_controller : component lab3_sopc_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => pll_c0_clk,                         --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component lab3_sopc_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component lab3_sopc_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => pll_c0_clk,                         --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	cpu_debug_reset_request_reset_ports_inv <= not cpu_debug_reset_request_reset;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_sdram_ctrl_s1_read_ports_inv <= not mm_interconnect_0_sdram_ctrl_s1_read;

	mm_interconnect_0_sdram_ctrl_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_ctrl_s1_byteenable;

	mm_interconnect_0_sdram_ctrl_s1_write_ports_inv <= not mm_interconnect_0_sdram_ctrl_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

end architecture rtl; -- of lab3_sopc
